`timescale 1ns / 1ps
module gelu_lut_module (
    input                       clk,
    input                       rst_n,
    input                       in_valid,     
    input      signed [15:0]    in_data,      
    output reg                  out_valid, 
    output reg signed [10:0]    out_data    
);

    //logic signed [15:0] gelu_rom [0:1280];
    localparam signed [10:0] gelu_rom [0:1279] = '{
    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFC,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFB,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFFA,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF9,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF7,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF6,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF5,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF3,    16'hFFF3,    16'hFFF3,    16'hFFF3,    16'hFFF3,    16'hFFF3,    16'hFFF3,    16'hFFF3,    16'hFFF3,    16'hFFF3,    16'hFFF3,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF1,    16'hFFF1,    16'hFFF1,    16'hFFF1,    16'hFFF1,    16'hFFF1,    16'hFFF1,    16'hFFF1,    16'hFFF1,    16'hFFF1,    16'hFFF0,    16'hFFF0,    16'hFFF0,    16'hFFF0,    16'hFFF0,    16'hFFF0,    16'hFFF0,    16'hFFF0,    16'hFFF0,    16'hFFEF,    16'hFFEF,    16'hFFEF,    16'hFFEF,    16'hFFEF,    16'hFFEF,    16'hFFEF,    16'hFFEF,    16'hFFEF,    16'hFFEE,    16'hFFEE,    16'hFFEE,    16'hFFEE,    16'hFFEE,    16'hFFEE,    16'hFFEE,    16'hFFEE,    16'hFFEE,    16'hFFED,    16'hFFED,    16'hFFED,    16'hFFED,    16'hFFED,    16'hFFED,    16'hFFED,    16'hFFED,    16'hFFED,    16'hFFEC,    16'hFFEC,    16'hFFEC,    16'hFFEC,    16'hFFEC,    16'hFFEC,    16'hFFEC,    16'hFFEC,    16'hFFEC,    16'hFFEB,    16'hFFEB,    16'hFFEB,    16'hFFEB,    16'hFFEB,    16'hFFEB,    16'hFFEB,    16'hFFEB,    16'hFFEA,    16'hFFEA,    16'hFFEA,    16'hFFEA,    16'hFFEA,    16'hFFEA,    16'hFFEA,    16'hFFEA,    16'hFFE9,    16'hFFE9,    16'hFFE9,    16'hFFE9,    16'hFFE9,    16'hFFE9,    16'hFFE9,    16'hFFE9,    16'hFFE8,    16'hFFE8,    16'hFFE8,    16'hFFE8,    16'hFFE8,    16'hFFE8,    16'hFFE8,    16'hFFE8,    16'hFFE7,    16'hFFE7,    16'hFFE7,    16'hFFE7,    16'hFFE7,    16'hFFE7,    16'hFFE7,    16'hFFE7,    16'hFFE6,    16'hFFE6,    16'hFFE6,    16'hFFE6,    16'hFFE6,    16'hFFE6,    16'hFFE6,    16'hFFE6,    16'hFFE5,    16'hFFE5,    16'hFFE5,    16'hFFE5,    16'hFFE5,    16'hFFE5,    16'hFFE5,    16'hFFE5,    16'hFFE4,    16'hFFE4,    16'hFFE4,    16'hFFE4,    16'hFFE4,    16'hFFE4,    16'hFFE4,    16'hFFE4,    16'hFFE3,    16'hFFE3,    16'hFFE3,    16'hFFE3,    16'hFFE3,    16'hFFE3,    16'hFFE3,    16'hFFE2,    16'hFFE2,    16'hFFE2,    16'hFFE2,    16'hFFE2,    16'hFFE2,    16'hFFE2,    16'hFFE2,    16'hFFE1,    16'hFFE1,    16'hFFE1,    16'hFFE1,    16'hFFE1,    16'hFFE1,    16'hFFE1,    16'hFFE1,    16'hFFE0,    16'hFFE0,    16'hFFE0,    16'hFFE0,    16'hFFE0,    16'hFFE0,    16'hFFE0,    16'hFFE0,    16'hFFDF,    16'hFFDF,    16'hFFDF,    16'hFFDF,    16'hFFDF,    16'hFFDF,    16'hFFDF,    16'hFFDF,    16'hFFDE,    16'hFFDE,    16'hFFDE,    16'hFFDE,    16'hFFDE,    16'hFFDE,    16'hFFDE,    16'hFFDE,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDC,    16'hFFDC,    16'hFFDC,    16'hFFDC,    16'hFFDC,    16'hFFDC,    16'hFFDC,    16'hFFDC,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD4,    16'hFFD4,    16'hFFD4,    16'hFFD4,    16'hFFD4,    16'hFFD4,    16'hFFD4,    16'hFFD4,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD5,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD6,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD7,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD8,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFD9,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDA,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDB,    16'hFFDC,    16'hFFDC,    16'hFFDC,    16'hFFDC,    16'hFFDC,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDD,    16'hFFDE,    16'hFFDE,    16'hFFDE,    16'hFFDE,    16'hFFDE,    16'hFFDF,    16'hFFDF,    16'hFFDF,    16'hFFDF,    16'hFFE0,    16'hFFE0,    16'hFFE0,    16'hFFE0,    16'hFFE1,    16'hFFE1,    16'hFFE1,    16'hFFE1,    16'hFFE2,    16'hFFE2,    16'hFFE2,    16'hFFE2,    16'hFFE3,    16'hFFE3,    16'hFFE3,    16'hFFE3,    16'hFFE4,    16'hFFE4,    16'hFFE4,    16'hFFE5,    16'hFFE5,    16'hFFE5,    16'hFFE5,    16'hFFE6,    16'hFFE6,    16'hFFE6,    16'hFFE7,    16'hFFE7,    16'hFFE7,    16'hFFE8,    16'hFFE8,    16'hFFE8,    16'hFFE9,    16'hFFE9,    16'hFFE9,    16'hFFEA,    16'hFFEA,    16'hFFEA,    16'hFFEB,    16'hFFEB,    16'hFFEB,    16'hFFEC,    16'hFFEC,    16'hFFEC,    16'hFFED,    16'hFFED,    16'hFFED,    16'hFFEE,    16'hFFEE,    16'hFFEE,    16'hFFEF,    16'hFFEF,    16'hFFF0,    16'hFFF0,    16'hFFF0,    16'hFFF1,    16'hFFF1,    16'hFFF2,    16'hFFF2,    16'hFFF2,    16'hFFF3,    16'hFFF3,    16'hFFF4,    16'hFFF4,    16'hFFF4,    16'hFFF5,    16'hFFF5,    16'hFFF6,    16'hFFF6,    16'hFFF7,    16'hFFF7,    16'hFFF8,    16'hFFF8,    16'hFFF8,    16'hFFF9,    16'hFFF9,    16'hFFFA,    16'hFFFA,    16'hFFFB,    16'hFFFB,    16'hFFFC,    16'hFFFC,    16'hFFFD,    16'hFFFD,    16'hFFFE,    16'hFFFE,    16'hFFFF,    16'hFFFF,    16'h0000,    16'h0000,    16'h0001,    16'h0001,    16'h0002,    16'h0002,    16'h0003,    16'h0003,    16'h0004,    16'h0004,    16'h0005,    16'h0005,    16'h0006,    16'h0006,    16'h0007,    16'h0007,    16'h0008,    16'h0008,    16'h0009,    16'h000A,    16'h000A,    16'h000B,    16'h000B,    16'h000C,    16'h000C,    16'h000D,    16'h000D,    16'h000E,    16'h000F,    16'h000F,    16'h0010,    16'h0010,    16'h0011,    16'h0012,    16'h0012,    16'h0013,    16'h0013,    16'h0014,    16'h0015,    16'h0015,    16'h0016,    16'h0016,    16'h0017,    16'h0018,    16'h0018,    16'h0019,    16'h001A,    16'h001A,    16'h001B,    16'h001C,    16'h001C,    16'h001D,    16'h001E,    16'h001E,    16'h001F,    16'h0020,    16'h0020,    16'h0021,    16'h0022,    16'h0022,    16'h0023,    16'h0024,    16'h0024,    16'h0025,    16'h0026,    16'h0026,    16'h0027,    16'h0028,    16'h0028,    16'h0029,    16'h002A,    16'h002B,    16'h002B,    16'h002C,    16'h002D,    16'h002D,    16'h002E,    16'h002F,    16'h0030,    16'h0030,    16'h0031,    16'h0032,    16'h0033,    16'h0033,    16'h0034,    16'h0035,    16'h0036,    16'h0036,    16'h0037,    16'h0038,    16'h0039,    16'h0039,    16'h003A,    16'h003B,    16'h003C,    16'h003C,    16'h003D,    16'h003E,    16'h003F,    16'h0040,    16'h0040,    16'h0041,    16'h0042,    16'h0043,    16'h0044,    16'h0044,    16'h0045,    16'h0046,    16'h0047,    16'h0048,    16'h0048,    16'h0049,    16'h004A,    16'h004B,    16'h004C,    16'h004D,    16'h004D,    16'h004E,    16'h004F,    16'h0050,    16'h0051,    16'h0052,    16'h0052,    16'h0053,    16'h0054,    16'h0055,    16'h0056,    16'h0057,    16'h0058,    16'h0059,    16'h0059,    16'h005A,    16'h005B,    16'h005C,    16'h005D,    16'h005E,    16'h005F,    16'h0060,    16'h0060,    16'h0061,    16'h0062,    16'h0063,    16'h0064,    16'h0065,    16'h0066,    16'h0067,    16'h0068,    16'h0069,    16'h0069,    16'h006A,    16'h006B,    16'h006C,    16'h006D,    16'h006E,    16'h006F,    16'h0070,    16'h0071,    16'h0072,    16'h0073,    16'h0074,    16'h0075,    16'h0075,    16'h0076,    16'h0077,    16'h0078,    16'h0079,    16'h007A,    16'h007B,    16'h007C,    16'h007D,    16'h007E,    16'h007F,    16'h0080,    16'h0081,    16'h0082,    16'h0083,    16'h0084,    16'h0085,    16'h0086,    16'h0087,    16'h0088,    16'h0089,    16'h008A,    16'h008B,    16'h008C,    16'h008D,    16'h008E,    16'h008F,    16'h0090,    16'h0091,    16'h0091,    16'h0092,    16'h0093,    16'h0094,    16'h0095,    16'h0096,    16'h0097,    16'h0098,    16'h009A,    16'h009B,    16'h009C,    16'h009D,    16'h009E,    16'h009F,    16'h00A0,    16'h00A1,    16'h00A2,    16'h00A3,    16'h00A4,    16'h00A5,    16'h00A6,    16'h00A7,    16'h00A8,    16'h00A9,    16'h00AA,    16'h00AB,    16'h00AC,    16'h00AD,    16'h00AE,    16'h00AF,    16'h00B0,    16'h00B1,    16'h00B2,    16'h00B3,    16'h00B4,    16'h00B5,    16'h00B6,    16'h00B7,    16'h00B8,    16'h00B9,    16'h00BB,    16'h00BC,    16'h00BD,    16'h00BE,    16'h00BF,    16'h00C0,    16'h00C1,    16'h00C2,    16'h00C3,    16'h00C4,    16'h00C5,    16'h00C6,    16'h00C7,    16'h00C8,    16'h00C9,    16'h00CA,    16'h00CC,    16'h00CD,    16'h00CE,    16'h00CF,    16'h00D0,    16'h00D1,    16'h00D2,    16'h00D3,    16'h00D4,    16'h00D5,    16'h00D6,    16'h00D7,    16'h00D8,    16'h00DA,    16'h00DB,    16'h00DC,    16'h00DD,    16'h00DE,    16'h00DF,    16'h00E0,    16'h00E1,    16'h00E2,    16'h00E3,    16'h00E4,    16'h00E6,    16'h00E7,    16'h00E8,    16'h00E9,    16'h00EA,    16'h00EB,    16'h00EC,    16'h00ED,    16'h00EE,    16'h00EF,    16'h00F1,    16'h00F2,    16'h00F3,    16'h00F4,    16'h00F5,    16'h00F6,    16'h00F7,    16'h00F8,    16'h00F9,    16'h00FA,    16'h00FC,    16'h00FD,    16'h00FE,    16'h00FF,    16'h0100,    16'h0101,    16'h0102,    16'h0103,    16'h0104,    16'h0106,    16'h0107,    16'h0108,    16'h0109,    16'h010A,    16'h010B,    16'h010C,    16'h010D,    16'h010F,    16'h0110,    16'h0111,    16'h0112,    16'h0113,    16'h0114,    16'h0115,    16'h0116,    16'h0117,    16'h0119,    16'h011A,    16'h011B,    16'h011C,    16'h011D,    16'h011E,    16'h011F,    16'h0120,    16'h0122,    16'h0123,    16'h0124,    16'h0125,    16'h0126,    16'h0127,    16'h0128,    16'h0129,    16'h012B,    16'h012C,    16'h012D,    16'h012E,    16'h012F,    16'h0130,    16'h0131,    16'h0132,    16'h0134,    16'h0135,    16'h0136,    16'h0137,    16'h0138,    16'h0139,    16'h013A,    16'h013B,    16'h013D,    16'h013E,    16'h013F,    16'h0140,    16'h0141,    16'h0142,    16'h0143,    16'h0144,    16'h0146,    16'h0147,    16'h0148,    16'h0149,    16'h014A,    16'h014B,    16'h014C,    16'h014E,    16'h014F,    16'h0150,    16'h0151,    16'h0152,    16'h0153,    16'h0154,    16'h0155,    16'h0157,    16'h0158,    16'h0159,    16'h015A,    16'h015B,    16'h015C,    16'h015D,    16'h015E,    16'h0160,    16'h0161,    16'h0162,    16'h0163,    16'h0164,    16'h0165,    16'h0166,    16'h0167,    16'h0169,    16'h016A,    16'h016B,    16'h016C,    16'h016D,    16'h016E,    16'h016F,    16'h0170,    16'h0172,    16'h0173,    16'h0174,    16'h0175,    16'h0176,    16'h0177,    16'h0178,    16'h0179,    16'h017B,    16'h017C,    16'h017D,    16'h017E,    16'h017F,    16'h0180,    16'h0181,    16'h0182,    16'h0184,    16'h0185,    16'h0186,    16'h0187,    16'h0188,    16'h0189,    16'h018A,    16'h018B,    16'h018D,    16'h018E,    16'h018F,    16'h0190,    16'h0191,    16'h0192,    16'h0193,    16'h0194,    16'h0196,    16'h0197,    16'h0198,    16'h0199,    16'h019A,    16'h019B,    16'h019C,    16'h019D,    16'h019E,    16'h01A0,    16'h01A1,    16'h01A2,    16'h01A3,    16'h01A4,    16'h01A5,    16'h01A6,    16'h01A7,    16'h01A8,    16'h01AA,    16'h01AB,    16'h01AC,    16'h01AD,    16'h01AE,    16'h01AF,    16'h01B0,    16'h01B1,    16'h01B2,    16'h01B4,    16'h01B5,    16'h01B6,    16'h01B7,    16'h01B8,    16'h01B9,    16'h01BA,    16'h01BB,    16'h01BC,    16'h01BE,    16'h01BF,    16'h01C0,    16'h01C1,    16'h01C2,    16'h01C3,    16'h01C4,    16'h01C5,    16'h01C6,    16'h01C8,    16'h01C9,    16'h01CA,    16'h01CB,    16'h01CC,    16'h01CD,    16'h01CE,    16'h01CF,    16'h01D0,    16'h01D1,    16'h01D3,    16'h01D4,    16'h01D5,    16'h01D6,    16'h01D7,    16'h01D8,    16'h01D9,    16'h01DA,    16'h01DB,    16'h01DC,    16'h01DD,    16'h01DF,    16'h01E0,    16'h01E1,    16'h01E2,    16'h01E3,    16'h01E4,    16'h01E5,    16'h01E6,    16'h01E7,    16'h01E8,    16'h01E9,    16'h01EB,    16'h01EC,    16'h01ED,    16'h01EE,    16'h01EF,    16'h01F0,    16'h01F1,    16'h01F2,    16'h01F3,    16'h01F4,    16'h01F5,    16'h01F7,    16'h01F8,    16'h01F9,    16'h01FA,    16'h01FB,    16'h01FC,    16'h01FD,    16'h01FE,    16'h01FF,    16'h0200,    16'h0201,    16'h0202,    16'h0204,    16'h0205,    16'h0206,    16'h0207,    16'h0208,    16'h0209,    16'h020A,    16'h020B,    16'h020C,    16'h020D,    16'h020E,    16'h020F,    16'h0210,    16'h0212,    16'h0213,    16'h0214,    16'h0215,    16'h0216,    16'h0217,    16'h0218,    16'h0219,    16'h021A,    16'h021B,    16'h021C,    16'h021D,    16'h021E,    16'h021F,    16'h0220,    16'h0222,    16'h0223,    16'h0224,    16'h0225,    16'h0226,    16'h0227,    16'h0228,    16'h0229,    16'h022A,    16'h022B,    16'h022C,    16'h022D,    16'h022E,    16'h022F,    16'h0230,    16'h0232,    16'h0233,    16'h0234,    16'h0235,    16'h0236,    16'h0237,    16'h0238,    16'h0239,    16'h023A,    16'h023B,    16'h023C,    16'h023D,    16'h023E,    16'h023F,    16'h0240,    16'h0241,    16'h0242,    16'h0244,    16'h0245,    16'h0246,    16'h0247,    16'h0248,    16'h0249,    16'h024A,    16'h024B,    16'h024C,    16'h024D,    16'h024E,    16'h024F,    16'h0250,    16'h0251,    16'h0252,    16'h0253,    16'h0254,    16'h0255,    16'h0256,    16'h0258,    16'h0259,    16'h025A,    16'h025B,    16'h025C,    16'h025D,    16'h025E,    16'h025F,    16'h0260,    16'h0261,    16'h0262,    16'h0263,    16'h0264,    16'h0265,    16'h0266,    16'h0267,    16'h0268,    16'h0269,    16'h026A,    16'h026B,    16'h026C,    16'h026D,    16'h026F,    16'h0270,    16'h0271,    16'h0272,    16'h0273,    16'h0274,    16'h0275,    16'h0276,    16'h0277,    16'h0278,    16'h0279,    16'h027A,    16'h027B};

    /*initial begin
        $readmemh("files/gelu_lut_hex_truncate.txt", gelu_rom);
    end*/
    // 將 in_data 轉換為 address
    // -32768 -> 0 
    // 0 -> 32768
    // 32767 -> 65535 
    logic [10:0] address_n, address;
    logic [15:0] out_data_n,out_valid_n;
    logic get_address, get_address_n;
    assign address_n = $unsigned(in_data) + 640;

    always_ff @(posedge clk,negedge rst_n) begin
        if(!rst_n)begin
            out_data<=0;
            out_valid<=0;
            address<=0;
            get_address<=0;
        end else begin
            out_data<=out_data_n;
            out_valid<=out_valid_n;
            address<=address_n;
            get_address<=get_address_n;
        end
    end
    always_comb begin 
        out_data_n = gelu_rom[address];
        get_address_n = 0;
        out_valid_n = 0;
        if(in_valid)begin
            get_address_n = 1;
        end
        if (get_address) begin
            out_valid_n = 1;
        end 
    end

endmodule